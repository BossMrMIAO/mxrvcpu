//********************************************************
// mxrv_ctrl
// function: decide when to send hold and flush command
//********************************************************


module mxrv_ctrl (
    ports
);
    
endmodule