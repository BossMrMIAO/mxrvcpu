
module axi_arbiter(
    input wire clk,
    input wire rst_n,
    input [31:0]    addr

);




endmodule