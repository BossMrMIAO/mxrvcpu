//********************************************************
// ctrl
// function: decide when to send hold and flush command
//********************************************************


module ctrl (

);
    
endmodule