//****************************************************
// if_id
// function:位于取指单元与译码单元之间，打一拍起到增加流水线级数作用
//****************************************************

module if_id #(
    
) (
    // global clock
    input clk,
    input rst_n,
    
);
    
endmodule